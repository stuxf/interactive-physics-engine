module main(
    // input logic SDI, SDO, SCLK, CE,
    output logic A, B, C, D, E,
    output logic R1, R2, B1, B2, G1, G2,
    output logic CLK, OE, LAT
);

endmodule
